module not_32bit(
	input [31:0] num,
	output [31:0] not_num);
	
	not(not_num[0],num[0]);
	not(not_num[1],num[1]);
	not(not_num[2],num[2]);
	not(not_num[3],num[3]);
	not(not_num[4],num[4]);
	not(not_num[5],num[5]);
	not(not_num[6],num[6]);
	not(not_num[7],num[7]);
	not(not_num[8],num[8]);
	not(not_num[9],num[9]);
	not(not_num[10],num[10]);
	not(not_num[11],num[11]);
	not(not_num[12],num[12]);
	not(not_num[13],num[13]);
	not(not_num[14],num[14]);
	not(not_num[15],num[15]);
	not(not_num[16],num[16]);
	not(not_num[17],num[17]);
	not(not_num[18],num[18]);
	not(not_num[19],num[19]);
	not(not_num[20],num[20]);
	not(not_num[21],num[21]);
	not(not_num[22],num[22]);
	not(not_num[23],num[23]);
	not(not_num[24],num[24]);
	not(not_num[25],num[25]);
	not(not_num[26],num[26]);
	not(not_num[27],num[27]);
	not(not_num[28],num[28]);
	not(not_num[29],num[29]);
	not(not_num[30],num[30]);
	not(not_num[31],num[31]);
	
endmodule
